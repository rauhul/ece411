module stage_writeback (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule