module xor2(
	input a, b,
	output f
);

assign f = a ^ b;

endmodule : xor2