module stage_execute (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule