module barrier_EX_MEM (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: barrier_EX_MEM