import lc3b_types::*;

module branch_predictor (
    /* INPUTS */

    /* OUTPUTS */
    output logic prediction
);

assign prediction = 0;

endmodule : branch_predictor
