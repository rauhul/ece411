module stage_decode (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule