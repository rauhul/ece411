module stage_ID (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: stage_ID