module stage_WB (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: stage_WB