module barrier_ID_EX (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: barrier_ID_EX