module barrier_IF_ID (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: barrier_IF_ID