module stage_mem (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule