module stage_EX (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: stage_EX