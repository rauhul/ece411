module barrier_MEM_WB (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: barrier_MEM_WB