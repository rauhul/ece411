module stage_IF (
    /* INPUTS */
    input clk

    /* OUTPUTS */
);

endmodule: stage_IF